module FP_acc(in1, in2, out);
parameter DATA_WIDTH = 32;
input 	[DATA_WIDTH-1:0] in1;// int_bits=4, frac_bits=28
input 	[DATA_WIDTH-1:0] in2;// single-precision floating-point
output reg [DATA_WIDTH-1:0] out;


always@(*) begin
	in1
end

endmodule